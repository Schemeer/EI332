library verilog;
use verilog.vl_types.all;
entity pipelined_computer_sim is
end pipelined_computer_sim;
