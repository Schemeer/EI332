library verilog;
use verilog.vl_types.all;
entity sc_computer_sim is
end sc_computer_sim;
